////////////////////////////////////////////////////////////////////////////////// Filename: man_dec.v// Description : Verilog module for Manchester code decoder// Author: LI Huang// Date: 4/29/2020////////////////////////////////////////////////////////////////////////////////`timescale 1ns/1psmodule man_dec(clk,rst,code,data,clk1);input   clk;    // clk from the internal oscillatorinput   rst;input   code;output  data;output  clk1;   // balanced data clkwire re_clk;    //recoverd clockwire o_reset;   //the final reset signalwire g_clk;     //gating clockwire [3:0]d_count;wire [3:0]c_count;wire d_comparison; wire c_comparison; reg dff1;reg [3:0]d_counter; //data counterreg [3:0]c_counter; //clock counterreg data_reg;reg clk1_reg;assign re_clk=data^code;assign g_clk=dff1&clk;assign d_comparison=(d_count>4'd12)? 0:1;  //data count comparatorassign c_comparison=(d_count>4'd8)? 0:1;  //balanced clock count comparatorassign o_reset=rst & d_comparison;//----------dff1 is the trigger of the data counter------// always @(posedge re_clk or negedge o_reset)    begin        if (!o_reset)            dff1<=0;        else            dff1<=1;    end//----------data conter------//always @(posedge g_clk or negedge o_reset)    begin        if (!o_reset)            d_counter<=0;        else            d_counter<=d_counter+1;    endassign d_count=d_counter;//----------data sampling register------//    always @(posedge d_comparison or negedge rst)    begin        if (!rst)            data_reg<= 0;        else            data_reg<=code;    endassign data=data_reg;    //----------balanced clock conter------//always @(posedge clk or posedge re_clk)    begin        if (re_clk)            c_counter<=0;        else             c_counter<=c_counter+1;    endassign c_count=c_counter;//----------balanced clock sampling register------//always @(posedge re_clk or negedge c_comparison)    begin        if(!c_comparison)            clk1_reg<=0;        else             clk1_reg<=1;    endassign clk1=clk1_reg;endmodule////////////////////////////////////////////////////////////////////////////////// Filename    : man_enc.v// Author      : lihuang       4/29/2020// Description : Verilog module for Manchester encoder////////////////////////////////////////////////////////////////////////////////`timescale 1ns/1psmodule man_enc (clk,rst,data,code);input clk;      //balanced clock from the decoderinput data;     //data from the decoder with matching phase with clkinput rst;output code;assign code=(!rst)? 0:             clk ~^ data;endmodule