////////////////////////////////////////////////////////////////////////////////// Filename : pwm_model.v// Author : lihuang 4//22/2020// Description : Verilog module for PMW wave forming////////////////////////////////////////////////////////////////////////////////
`timescale 1ns/1ns
module pwm_model(clk,rst,intensity,ctl);input clk;input rst;input [9:0]intensity;wire rst_2;wire [9:0]count;wire [15:0]inten_n;wire [15:0] sum;wire a;assign inten_n = ~ intensity;assign a=sum[10];//use asynchronized_reset and synchronized release to improve the robustnessarest_srls a1(.clk(clk),.rst(rst),.a(rst_2));//use the counter to count the value of input clock cyclescounter counter1(.clk(clk),.rst(rst_2),.count(count));//use the cla_16bit to form a sub which can perform the comparisoncla_16bit sub(.a(count),.b(inten_n),.cin(1),.sum(sum),.cout(),.pg(),.gg());//use the multiplexer to define the output signalmultipexer mul1(.a(a),.b(ctl));Endmodule////////////////////////////////////////////////////////////////////////////////// Filename : pwm.v// Author : lihuang 4/22/2020// Description : Verilog module for multiplexer////////////////////////////////////////////////////////////////////////////////module multipexer(a,b);input a;output b;assign b=(a==0)? 0:1;endmodule////////////////////////////////////////////////////////////////////////////////// Filename : arest_sls.v// Author : lihuang 4/22/2020// Description : Verilog module for asychronize reseting and sychronized releasing////////////////////////////////////////////////////////////////////////////////module arest_srls(clk,rst,a);input clk;input rst;output a;reg rst_1;reg rst_2; assign a = rst_2;always @(posedge clk or negedge rst)beginif (!rst)beginrst_1<=0;rst_2<=0;endelsebeginrst_1<=1;rst_2<=rst_1;endendendmodule////////////////////////////////////////////////////////////////////////////////// Filename : counter.v// Author : lihuang 4/22/2020// Description : Verilog module for counter////////////////////////////////////////////////////////////////////////////////module counter(clk,rst,count);input clk;input rst;output [9:0]count;reg [9:0]counter;wire rst_2;assign rst_2 = rst;assign count =counter;//use counter to define the period value of outputalways @ (posedge clk or negedge rst_2)beginif (!rst_2)begincounter<=0;endelse if (counter == {10{1'b1}}-1'b1)begincounter<=0;endelsebegincounter<=counter+1;endendendmodule////////////////////////////////////////////////////////////////////////////////// Filename : cla_16bit.v// Author : lihuang 4/22/2020// Description : Verilog module for cla_16bit////////////////////////////////////////////////////////////////////////////////module cla_16bit (a, b, cin, sum, cout, pg, gg);input [15:0] a;input [15:0] b;input cin;output [15:0] sum;output cout;output pg; //16-bit block group propagateoutput gg; //16-bit block group generatewire [3:0] p;wire [3:0] g;wire [4:0] c;assign cout=c[4];assign c[0]=cin;assign pg = &p;assign gg = g[3] | (g[2]&p[3]) | (g[1]&p[3]&p[2]) | (g[0]&p[3]&p[2]&p[1]);assign c[1] = g[0] | (p[0]&c[0]);assign c[2] = g[1] | (p[1]&g[0]) | (p[1]&p[0]&c[0]);assign c[3] = g[2] | (p[2]&g[1]) | (p[2]&p[1]&g[0]) | (p[2]&p[1]&p[0]&c[0]);assign c[4] = g[3] | (p[3]&g[2]) | (p[3]&p[2]&g[1]) | (p[3]&p[2]&p[1]&g[0])| (p[3]&p[2]&p[1]&p[0]&c[0]);cla_4bit cla0(.a(a[3:0]),.b(b[3:0]),.cin(c[0]),.sum(sum[3:0]),.cout(),.pg(p[0]),.gg(g[0]));cla_4bit cla1(.a(a[7:4]),.b(b[7:4]),.cin(c[1]),.sum(sum[7:4]),.cout(),.pg(p[1]),.gg(g[1]));cla_4bit cla2(.a(a[11:8]),.b(b[11:8]),.cin(c[2]),.sum(sum[11:8]),.cout(),.pg(p[2]),.gg(g[2]));cla_4bit cla3(.a(a[15:12]),.b(b[15:12]),.cin(c[3]),.sum(sum[15:12]),.cout(),.pg(p[3]),.gg(g[3]));Endmodule//------------4-bit CLA adder------------////------------the main advantage of CLA architecture is the reduction in carry generation time------------//module cla_4bit(a,b, cin, sum, cout, pg, gg);input [3:0] a;input [3:0] b;input cin;output [3:0] sum;output cout;output pg; //4-bit block group propagateoutput gg; //4-bit block group generatewire [3:0] p;wire [3:0] g;wire [4:0] c;//-----------stage1-----------////------------calculate generate and propagate in the same time-----------//assign p=a^b;assign g=a&b;assign sum = p[3:0]^c[3:0];assign cout=c[4];assign c[0]=cin;assign pg = &p;assign gg = g[3] | (g[2]&p[3]) | (g[1]&p[3]&p[2]) | (g[0]&p[3]&p[2]&p[1]);assign c[1] = g[0] | (p[0]&c[0]);assign c[2] = g[1] | (p[1]&g[0]) | (p[1]&p[0]&c[0]);assign c[3] = g[2] | (p[2]&g[1]) | (p[2]&p[1]&g[0]) | (p[2]&p[1]&p[0]&c[0]);assign c[4] = g[3] | (p[3]&g[2]) | (p[3]&p[2]&g[1]) | (p[3]&p[2]&p[1]&g[0]) | (p[3]&p[2]&p[1]&p[0]&c[0]);endmodule